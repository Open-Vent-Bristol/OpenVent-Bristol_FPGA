

library ieee;
use ieee.std_logic_1164.all;

ENTITY lps25h_baro_spi_format_tb IS
end entity lps25h_baro_spi_format_tb;


ARCHITECTURE testbench OF lps25h_baro_spi_format_tb IS
	constant MAX_DELAY: time := 100 ns;
	signal mstrclk: std_logic := '0';
	signal RST_L: std_logic := '0';
	signal BARO_OUT: std_logic := '0';
	signal baro_intr: std_logic := '0';
	signal	BARO_din: STD_LOGIC;
	signal	BARO_din_exp: STD_LOGIC;
	signal	BARO_SERCLK: STD_LOGIC;
	signal	BARO_SERCLK_exp: STD_LOGIC;
	signal	baro_CSN: STD_LOGIC;
	signal	baro_CSN_exp: STD_LOGIC;
	signal Press : STD_LOGIC_VECTOR(23 downto 0);
	signal Temp : STD_LOGIC_VECTOR(15 downto 0);
	signal AbsPress : STD_LOGIC_VECTOR(17 downto 0);

begin

--DUV instantiation
duv: entity work.LPS25H_BARO_spi_format port map(rst_L,mstrclk, baro_out, baro_INTR,baro_din, baro_serclk, baro_CSN, PRESS,TEMP,AbsPress);

--Stimuli generator
mstrclk <= not mstrclk after 100 ns;
RST_L <= '1' after 150 ns;
baro_INTR <=  '1' after	163	us,
'0' after	163.6	us, '1' after	740	us,
'0' after	748	us, '1' after	6803.6	us,
'0' after	6803.8	us, '1' after	7083	us,
'0' after	7087	us, '1' after	7333	us,
'0' after	7336	us;		

BARO_OUT <=  '1' after	165.5	us,
'0' after	167	us, '1' after	167.5	us,
'0' after	168	us, '1' after	168.5	us,
'0' after	169	us, '1' after	169.5	us,
'0' after	170	us, '1' after	170.5	us,
'0' after	171	us, '1' after	171.5	us,
'0' after	172	us, '1' after	172.5	us,
'0' after	173	us, '1' after	173.5	us,
'0' after	174	us, '1' after	174.5	us,
'0' after	175	us, '1' after	175.5	us,
'0' after	176	us, '1' after	176.5	us,
'0' after	177	us, '1' after	177.5	us,
'0' after	178	us, '1' after	178.5	us,
'0' after	179	us, '1' after	179.5	us,
'0' after	180	us, '1' after	180.5	us,
'0' after	181	us, '1' after	181.5	us,
'0' after	182	us, '1' after	182.5	us,
'0' after	183	us, '1' after	183.5	us,
'0' after	184	us, '1' after	184.5	us,
'0' after	185	us, '1' after	185.5	us,
'0' after	186	us, '1' after	186.5	us,
'0' after	187	us, '1' after	187.5	us,
'0' after	188	us, '1' after	188.5	us,
'0' after	189	us, '1' after	189.5	us,
'0' after	190	us, '1' after	190.5	us,
'0' after	191	us, '1' after	191.5	us,
'0' after	192	us, '1' after	192.5	us,
'0' after	193	us, '1' after	193.5	us,
'0' after	194	us, '1' after	194.5	us,
'0' after	195	us, '1' after	195.5	us,
'0' after	196	us, '1' after	196.5	us,
'0' after	197	us, '1' after	197.5	us,
'0' after	198	us, '1' after	198.5	us,
'0' after	199	us, '1' after	199.5	us,
'0' after	200	us, '1' after	200.5	us,
'0' after	201	us, '1' after	201.5	us,
'0' after	202	us, '1' after	202.5	us,
'0' after	203	us, '1' after	203.5	us,
'0' after	204	us, '1' after	204.5	us,
'0' after	205	us, '1' after	205.5	us,
'0' after	206	us, '1' after	206.5	us,
'0' after	207	us, '1' after	207.5	us,
'0' after	208	us, '1' after	208.5	us,
'0' after	209	us, '1' after	209.5	us,
'0' after	210	us, '1' after	210.5	us,
'0' after	211	us, '1' after	211.5	us,
'0' after	212	us, '1' after	212.5	us,
'0' after	213	us, '1' after	213.5	us,
'0' after	214	us, '1' after	214.5	us,
'0' after	215	us, '1' after	215.5	us,
'0' after	216	us, '1' after	216.5	us,
'0' after	217	us, '1' after	217.5	us,
'0' after	218	us, '1' after	218.5	us,
'0' after	219	us, '1' after	219.5	us,
'0' after	220	us, '1' after	220.5	us,
'0' after	221	us, '1' after	221.5	us,
'0' after	222	us, '1' after	222.5	us,
'0' after	223	us, '1' after	223.5	us,
'0' after	224	us, '1' after	224.5	us,
'0' after	225	us, '1' after	225.5	us,
'0' after	226	us, '1' after	226.5	us,
'0' after	227	us, '1' after	227.5	us,
'0' after	228	us, '1' after	228.5	us,
'0' after	229	us, '1' after	229.5	us,
'0' after	230	us, '1' after	230.5	us,
'0' after	231	us, '1' after	231.5	us,
'0' after	232	us, '1' after	232.5	us,
'0' after	233	us, '1' after	233.5	us,
'0' after	234	us, '1' after	234.5	us,
'0' after	235	us, '1' after	235.5	us,
'0' after	236	us, '1' after	236.5	us,
'0' after	237	us, '1' after	237.5	us,
'0' after	238	us, '1' after	238.5	us,
'0' after	239	us, '1' after	239.5	us,
'0' after	240	us, '1' after	240.5	us,
'0' after	241	us, '1' after	241.5	us,
'0' after	242	us, '1' after	242.5	us,
'0' after	243	us, '1' after	243.5	us,
'0' after	244	us, '1' after	244.5	us,
'0' after	245	us, '1' after	245.5	us,
'0' after	246	us, '1' after	246.5	us,
'0' after	247	us, '1' after	247.5	us,
'0' after	248	us, '1' after	248.5	us,
'0' after	249	us, '1' after	249.5	us,
'0' after	250	us, '1' after	250.5	us,
'0' after	251	us, '1' after	251.5	us,
'0' after	252	us, '1' after	742.5	us,
'0' after	743	us, '1' after	743.5	us,
'0' after	744	us, '1' after	744.5	us,
'0' after	745	us, '1' after	745.5	us,
'0' after	746	us, '1' after	746.5	us,
'0' after	747	us, '1' after	747.5	us,
'0' after	748	us, '1' after	748.5	us,
'0' after	749	us, '1' after	749.5	us,
'0' after	750	us, '1' after	750.5	us,
'0' after	751	us, '1' after	751.5	us,
'0' after	752	us, '1' after	752.5	us,
'0' after	753	us, '1' after	753.5	us,
'0' after	754	us, '1' after	754.5	us,
'0' after	755	us, '1' after	755.5	us,
'0' after	756	us, '1' after	756.5	us,
'0' after	757	us, '1' after	757.5	us,
'0' after	758	us, '1' after	758.5	us,
'0' after	759	us, '1' after	759.5	us,
'0' after	760	us, '1' after	760.5	us,
'0' after	761	us, '1' after	761.5	us,
'0' after	762	us, '1' after	762.5	us,
'0' after	763	us, '1' after	763.5	us,
'0' after	764	us, '1' after	764.5	us,
'0' after	765	us, '1' after	765.5	us,
'0' after	766	us, '1' after	766.5	us,
'0' after	767	us, '1' after	767.5	us,
'0' after	768	us, '1' after	768.5	us,
'0' after	769	us, '1' after	769.5	us,
'0' after	770	us, '1' after	770.5	us,
'0' after	771	us, '1' after	771.5	us,
'0' after	772	us, '1' after	772.5	us,
'0' after	773	us, '1' after	773.5	us,
'0' after	774	us, '1' after	774.5	us,
'0' after	775	us, '1' after	775.5	us,
'0' after	776	us, '1' after	776.5	us,
'0' after	777	us, '1' after	777.5	us,
'0' after	778	us, '1' after	778.5	us,
'0' after	779	us, '1' after	779.5	us,
'0' after	780	us, '1' after	780.5	us,
'0' after	781	us, '1' after	781.5	us,
'0' after	782	us, '1' after	782.5	us,
'0' after	783	us, '1' after	783.5	us,
'0' after	784	us, '1' after	784.5	us,
'0' after	785	us, '1' after	785.5	us,
'0' after	786	us, '1' after	786.5	us,
'0' after	787	us, '1' after	787.5	us,
'0' after	788	us, '1' after	788.5	us,
'0' after	789	us, '1' after	789.5	us,
'0' after	790	us, '1' after	790.5	us,
'0' after	791	us, '1' after	791.5	us,
'0' after	792	us, '1' after	792.5	us,
'0' after	793	us, '1' after	793.5	us,
'0' after	794	us, '1' after	794.5	us,
'0' after	795	us, '1' after	795.5	us,
'0' after	796	us, '1' after	796.5	us,
'0' after	797	us, '1' after	797.5	us,
'0' after	798	us, '1' after	798.5	us,
'0' after	799	us, '1' after	799.5	us,
'0' after	800	us, '1' after	800.5	us,
'0' after	801	us, '1' after	801.5	us,
'0' after	802	us, '1' after	802.5	us,
'0' after	803	us, '1' after	803.5	us,
'0' after	804	us, '1' after	804.5	us,
'0' after	805	us, '1' after	805.5	us,
'0' after	806	us, '1' after	806.5	us,
'0' after	807	us, '1' after	807.5	us,
'0' after	808	us, '1' after	808.5	us,
'0' after	809	us, '1' after	809.5	us,
'0' after	810	us, '1' after	810.5	us,
'0' after	811	us, '1' after	811.5	us,
'0' after	812	us, '1' after	812.5	us,
'0' after	813	us, '1' after	813.5	us,
'0' after	814	us, '1' after	814.5	us,
'0' after	815	us, '1' after	815.5	us,
'0' after	816	us, '1' after	816.5	us,
'0' after	817	us, '1' after	817.5	us,
'0' after	818	us, '1' after	818.5	us,
'0' after	819	us, '1' after	819.5	us,
'0' after	820	us, '1' after	820.5	us,
'0' after	821	us, '1' after	821.5	us,
'0' after	822	us, '1' after	822.5	us,
'0' after	823	us, '1' after	823.5	us,
'0' after	824	us, '1' after	824.5	us,
'0' after	825	us, '1' after	825.5	us,
'0' after	826	us, '1' after	826.5	us,
'0' after	827	us, '1' after	827.5	us,
'0' after	828	us, '1' after	828.5	us,
'0' after	829	us, '1' after	829.5	us,
'0' after	830	us, '1' after	6806.5	us,
'0' after	6807	us, '1' after	6807.5	us,
'0' after	6808	us, '1' after	6808.5	us,
'0' after	6809	us, '1' after	6809.5	us,
'0' after	6810	us, '1' after	6810.5	us,
'0' after	6811	us, '1' after	6811.5	us,
'0' after	6812	us, '1' after	6812.5	us,
'0' after	6813	us, '1' after	6813.5	us,
'0' after	6814	us, '1' after	6814.5	us,
'0' after	6815	us, '1' after	6815.5	us,
'0' after	6816	us, '1' after	6816.5	us,
'0' after	6817	us, '1' after	6817.5	us,
'0' after	6818	us, '1' after	6818.5	us,
'0' after	6819	us, '1' after	6819.5	us,
'0' after	6820	us, '1' after	6820.5	us,
'0' after	6821	us, '1' after	6821.5	us,
'0' after	6822	us, '1' after	6822.5	us,
'0' after	6823	us, '1' after	6823.5	us,
'0' after	6824	us, '1' after	6824.5	us,
'0' after	6825	us, '1' after	6825.5	us,
'0' after	6826	us, '1' after	6826.5	us,
'0' after	6827	us, '1' after	6827.5	us,
'0' after	6828	us, '1' after	6828.5	us,
'0' after	6829	us, '1' after	6829.5	us,
'0' after	6830	us, '1' after	6830.5	us,
'0' after	6831	us, '1' after	6831.5	us,
'0' after	6832	us, '1' after	6832.5	us,
'0' after	6833	us, '1' after	6833.5	us,
'0' after	6834	us, '1' after	6834.5	us,
'0' after	6835	us, '1' after	6835.5	us,
'0' after	6836	us, '1' after	6836.5	us,
'0' after	6837	us, '1' after	6837.5	us,
'0' after	6838	us, '1' after	6838.5	us,
'0' after	6839	us, '1' after	6839.5	us,
'0' after	6840	us, '1' after	6840.5	us,
'0' after	6841	us, '1' after	6841.5	us,
'0' after	6842	us, '1' after	6842.5	us,
'0' after	6843	us, '1' after	6843.5	us,
'0' after	6844	us, '1' after	6844.5	us,
'0' after	6845	us, '1' after	6845.5	us,
'0' after	6846	us, '1' after	6846.5	us,
'0' after	6847	us, '1' after	6847.5	us,
'0' after	6848	us, '1' after	6848.5	us,
'0' after	6849	us, '1' after	6849.5	us,
'0' after	6850	us, '1' after	6850.5	us,
'0' after	6851	us, '1' after	6851.5	us,
'0' after	6852	us, '1' after	6852.5	us,
'0' after	6853	us, '1' after	6853.5	us,
'0' after	6854	us, '1' after	6854.5	us,
'0' after	6855	us, '1' after	6855.5	us,
'0' after	6856	us, '1' after	6856.5	us,
'0' after	6857	us, '1' after	6857.5	us,
'0' after	6858	us, '1' after	6858.5	us,
'0' after	6859	us, '1' after	6859.5	us,
'0' after	6860	us, '1' after	6860.5	us,
'0' after	6861	us, '1' after	6861.5	us,
'0' after	6862	us, '1' after	6862.5	us,
'0' after	6863	us, '1' after	6863.5	us,
'0' after	6864	us, '1' after	6864.5	us,
'0' after	6865	us, '1' after	6865.5	us,
'0' after	6866	us, '1' after	6866.5	us,
'0' after	6867	us, '1' after	6867.5	us,
'0' after	6868	us, '1' after	6868.5	us,
'0' after	6869	us, '1' after	6869.5	us,
'0' after	6870	us, '1' after	6870.5	us,
'0' after	6871	us, '1' after	6871.5	us,
'0' after	6872	us, '1' after	6872.5	us,
'0' after	6873	us, '1' after	6873.5	us,
'0' after	6874	us, '1' after	6874.5	us,
'0' after	6875	us, '1' after	6875.5	us,
'0' after	6876	us, '1' after	6876.5	us,
'0' after	6877	us, '1' after	6877.5	us,
'0' after	6878	us, '1' after	6878.5	us,
'0' after	6879	us, '1' after	6879.5	us,
'0' after	6880	us, '1' after	6880.5	us,
'0' after	6881	us, '1' after	6881.5	us,
'0' after	6882	us, '1' after	6882.5	us,
'0' after	6883	us, '1' after	6883.5	us,
'0' after	6884	us, '1' after	6884.5	us,
'0' after	6885	us, '1' after	6885.5	us,
'0' after	6886	us, '1' after	6886.5	us,
'0' after	6887	us, '1' after	6887.5	us,
'0' after	6888	us, '1' after	6888.5	us,
'0' after	6889	us, '1' after	6889.5	us,
'0' after	6890	us, '1' after	6890.5	us,
'0' after	6891	us, '1' after	6891.5	us,
'0' after	6892	us, '1' after	6892.5	us,
'0' after	6893	us, '1' after	7085.5	us,
'0' after	7086	us, '1' after	7086.5	us,
'0' after	7087	us, '1' after	7087.5	us,
'0' after	7088	us, '1' after	7088.5	us,
'0' after	7089	us, '1' after	7089.5	us,
'0' after	7090	us, '1' after	7090.5	us,
'0' after	7091	us, '1' after	7091.5	us,
'0' after	7092	us, '1' after	7092.5	us,
'0' after	7093	us, '1' after	7093.5	us,
'0' after	7094	us, '1' after	7094.5	us,
'0' after	7095	us, '1' after	7095.5	us,
'0' after	7096	us, '1' after	7096.5	us,
'0' after	7097	us, '1' after	7097.5	us,
'0' after	7098	us, '1' after	7098.5	us,
'0' after	7099	us, '1' after	7099.5	us,
'0' after	7100	us, '1' after	7100.5	us,
'0' after	7101	us, '1' after	7101.5	us,
'0' after	7102	us, '1' after	7102.5	us,
'0' after	7103	us, '1' after	7103.5	us,
'0' after	7104	us, '1' after	7104.5	us,
'0' after	7105	us, '1' after	7105.5	us,
'0' after	7106	us, '1' after	7106.5	us,
'0' after	7107	us, '1' after	7107.5	us,
'0' after	7108	us, '1' after	7108.5	us,
'0' after	7109	us, '1' after	7109.5	us,
'0' after	7110	us, '1' after	7110.5	us,
'0' after	7111	us, '1' after	7111.5	us,
'0' after	7112	us, '1' after	7112.5	us,
'0' after	7113	us, '1' after	7113.5	us,
'0' after	7114	us, '1' after	7114.5	us,
'0' after	7115	us, '1' after	7115.5	us,
'0' after	7116	us, '1' after	7116.5	us,
'0' after	7117	us, '1' after	7117.5	us,
'0' after	7118	us, '1' after	7118.5	us,
'0' after	7119	us, '1' after	7119.5	us,
'0' after	7120	us, '1' after	7120.5	us,
'0' after	7121	us, '1' after	7121.5	us,
'0' after	7122	us, '1' after	7122.5	us,
'0' after	7123	us, '1' after	7123.5	us,
'0' after	7124	us, '1' after	7124.5	us,
'0' after	7125	us, '1' after	7125.5	us,
'0' after	7126	us, '1' after	7126.5	us,
'0' after	7127	us, '1' after	7127.5	us,
'0' after	7128	us, '1' after	7128.5	us,
'0' after	7129	us, '1' after	7129.5	us,
'0' after	7130	us, '1' after	7130.5	us,
'0' after	7131	us, '1' after	7131.5	us,
'0' after	7132	us, '1' after	7132.5	us,
'0' after	7133	us, '1' after	7133.5	us,
'0' after	7134	us, '1' after	7134.5	us,
'0' after	7135	us, '1' after	7135.5	us,
'0' after	7136	us, '1' after	7136.5	us,
'0' after	7137	us, '1' after	7137.5	us,
'0' after	7138	us, '1' after	7138.5	us,
'0' after	7139	us, '1' after	7139.5	us,
'0' after	7140	us, '1' after	7140.5	us,
'0' after	7141	us, '1' after	7141.5	us,
'0' after	7142	us, '1' after	7142.5	us,
'0' after	7143	us, '1' after	7143.5	us,
'0' after	7144	us, '1' after	7144.5	us,
'0' after	7145	us, '1' after	7145.5	us,
'0' after	7146	us, '1' after	7146.5	us,
'0' after	7147	us, '1' after	7147.5	us,
'0' after	7148	us, '1' after	7148.5	us,
'0' after	7149	us, '1' after	7149.5	us,
'0' after	7150	us, '1' after	7150.5	us,
'0' after	7151	us, '1' after	7151.5	us,
'0' after	7152	us, '1' after	7152.5	us,
'0' after	7153	us, '1' after	7153.5	us,
'0' after	7154	us, '1' after	7154.5	us,
'0' after	7155	us, '1' after	7155.5	us,
'0' after	7156	us, '1' after	7156.5	us,
'0' after	7157	us, '1' after	7157.5	us,
'0' after	7158	us, '1' after	7158.5	us,
'0' after	7159	us, '1' after	7159.5	us,
'0' after	7160	us, '1' after	7160.5	us,
'0' after	7161	us, '1' after	7161.5	us,
'0' after	7162	us, '1' after	7162.5	us,
'0' after	7163	us, '1' after	7163.5	us,
'0' after	7164	us, '1' after	7164.5	us,
'0' after	7165	us, '1' after	7165.5	us,
'0' after	7166	us, '1' after	7166.5	us,
'0' after	7167	us, '1' after	7167.5	us,
'0' after	7168	us, '1' after	7168.5	us,
'0' after	7169	us, '1' after	7169.5	us,
'0' after	7170	us, '1' after	7170.5	us,
'0' after	7171	us, '1' after	7171.5	us,
'0' after	7172	us, '1' after	7335.5	us,
'0' after	7336	us, '1' after	7336.5	us,
'0' after	7337	us, '1' after	7337.5	us,
'0' after	7338	us, '1' after	7338.5	us,
'0' after	7339	us, '1' after	7339.5	us,
'0' after	7340	us, '1' after	7340.5	us,
'0' after	7341	us, '1' after	7341.5	us,
'0' after	7342	us, '1' after	7342.5	us,
'0' after	7343	us, '1' after	7343.5	us,
'0' after	7344	us, '1' after	7344.5	us,
'0' after	7345	us, '1' after	7345.5	us,
'0' after	7346	us, '1' after	7346.5	us,
'0' after	7347	us, '1' after	7347.5	us,
'0' after	7348	us, '1' after	7348.5	us,
'0' after	7349	us, '1' after	7349.5	us,
'0' after	7350	us, '1' after	7350.5	us,
'0' after	7351	us, '1' after	7351.5	us,
'0' after	7352	us, '1' after	7352.5	us,
'0' after	7353	us, '1' after	7353.5	us,
'0' after	7354	us, '1' after	7354.5	us,
'0' after	7355	us, '1' after	7355.5	us,
'0' after	7356	us, '1' after	7356.5	us,
'0' after	7357	us, '1' after	7357.5	us,
'0' after	7358	us, '1' after	7358.5	us,
'0' after	7359	us, '1' after	7359.5	us,
'0' after	7360	us, '1' after	7360.5	us,
'0' after	7361	us, '1' after	7361.5	us,
'0' after	7362	us, '1' after	7362.5	us,
'0' after	7363	us, '1' after	7363.5	us,
'0' after	7364	us, '1' after	7364.5	us,
'0' after	7365	us, '1' after	7365.5	us,
'0' after	7366	us, '1' after	7366.5	us,
'0' after	7367	us, '1' after	7367.5	us,
'0' after	7368	us, '1' after	7368.5	us,
'0' after	7369	us, '1' after	7369.5	us,
'0' after	7370	us, '1' after	7370.5	us,
'0' after	7371	us, '1' after	7371.5	us,
'0' after	7372	us, '1' after	7372.5	us,
'0' after	7373	us, '1' after	7373.5	us,
'0' after	7374	us, '1' after	7374.5	us,
'0' after	7375	us, '1' after	7375.5	us,
'0' after	7376	us, '1' after	7376.5	us,
'0' after	7377	us, '1' after	7377.5	us,
'0' after	7378	us, '1' after	7378.5	us,
'0' after	7379	us, '1' after	7379.5	us,
'0' after	7380	us, '1' after	7380.5	us,
'0' after	7381	us, '1' after	7381.5	us,
'0' after	7382	us, '1' after	7382.5	us,
'0' after	7383	us, '1' after	7383.5	us,
'0' after	7384	us, '1' after	7384.5	us,
'0' after	7385	us, '1' after	7385.5	us,
'0' after	7386	us, '1' after	7386.5	us,
'0' after	7387	us, '1' after	7387.5	us,
'0' after	7388	us, '1' after	7388.5	us,
'0' after	7389	us, '1' after	7389.5	us,
'0' after	7390	us, '1' after	7390.5	us,
'0' after	7391	us, '1' after	7391.5	us,
'0' after	7392	us, '1' after	7392.5	us,
'0' after	7393	us, '1' after	7393.5	us,
'0' after	7394	us, '1' after	7394.5	us,
'0' after	7395	us, '1' after	7395.5	us,
'0' after	7396	us, '1' after	7396.5	us,
'0' after	7397	us, '1' after	7397.5	us,
'0' after	7398	us, '1' after	7398.5	us,
'0' after	7399	us, '1' after	7399.5	us,
'0' after	7400	us, '1' after	7400.5	us,
'0' after	7401	us, '1' after	7401.5	us,
'0' after	7402	us, '1' after	7402.5	us,
'0' after	7403	us, '1' after	7403.5	us,
'0' after	7404	us, '1' after	7404.5	us,
'0' after	7405	us, '1' after	7405.5	us,
'0' after	7406	us, '1' after	7406.5	us,
'0' after	7407	us, '1' after	7407.5	us,
'0' after	7408	us, '1' after	7408.5	us,
'0' after	7409	us, '1' after	7409.5	us,
'0' after	7410	us, '1' after	7410.5	us,
'0' after	7411	us, '1' after	7411.5	us,
'0' after	7412	us, '1' after	7412.5	us,
'0' after	7413	us, '1' after	7413.5	us,
'0' after	7414	us, '1' after	7414.5	us,
'0' after	7415	us, '1' after	7415.5	us,
'0' after	7416	us, '1' after	7416.5	us,
'0' after	7417	us, '1' after	7417.5	us,
'0' after	7418	us, '1' after	7418.5	us,
'0' after	7419	us, '1' after	7419.5	us,
'0' after	7420	us, '1' after	7420.5	us,
'0' after	7421	us, '1' after	7421.5	us,
'0' after	7422	US;		

--Template Generator
BARO_DIN_exp <=  '1' after	4	us,
'0' after	5.3	us, '1' after	8	us,
'0' after	10.1	us, '1' after	23.2	us,
'0' after	24.5	us, '1' after	30.4	us,
'0' after	34.1	us, '1' after	40.8	us,
'0' after	42.1	us, '1' after	49.6	us,
'0' after	50.9	us, '1' after	59.2	us,
'0' after	60.5	us, '1' after	63.2	us,
'0' after	66.9	us, '1' after	77.6	us,
'0' after	78.9	us, '1' after	80.8	us,
'0' after	82.1	us, '1' after	82.4	us,
'0' after	83.7	us, '1' after	96	us,
'0' after	97.3	us, '1' after	99.2	us,
'0' after	101.3	us, '1' after	106.4	us,
'0' after	107.7	us, '1' after	114.4	us,
'0' after	115.7	us, '1' after	116.8	us,
'0' after	118.1	us, '1' after	132.8	us,
'0' after	134.1	us, '1' after	134.4	us,
'0' after	137.3	us, '1' after	137.6	us,
'0' after	139.7	us, '1' after	140	us,
'0' after	144.5	us, '1' after	165.6	us,
'0' after	166.9	us, '1' after	167.2	us,
'0' after	168.5	us, '1' after	168.8	us,
'0' after	170.1	us, '1' after	184	us,
'0' after	185.3	us, '1' after	185.6	us,
'0' after	186.9	us, '1' after	187.2	us,
'0' after	188.5	us, '1' after	189.6	us,
'0' after	190.9	us, '1' after	202.4	us,
'0' after	203.7	us, '1' after	204	us,
'0' after	205.3	us, '1' after	205.6	us,
'0' after	206.9	us, '1' after	207.2	us,
'0' after	208.5	us, '1' after	220.8	us,
'0' after	222.1	us, '1' after	222.4	us,
'0' after	223.7	us, '1' after	224	us,
'0' after	225.3	us, '1' after	225.6	us,
'0' after	227.7	us, '1' after	239.2	us,
'0' after	240.5	us, '1' after	240.8	us,
'0' after	242.1	us, '1' after	242.4	us,
'0' after	244.5	us, '1' after	742.4	us,
'0' after	743.7	us, '1' after	744	us,
'0' after	745.3	us, '1' after	745.6	us,
'0' after	746.9	us, '1' after	760.8	us,
'0' after	762.1	us, '1' after	762.4	us,
'0' after	763.7	us, '1' after	764	us,
'0' after	764.3	us, '1' after	766.4	us,
'0' after	767.7	us, '1' after	779.2	us,
'0' after	780.5	us, '1' after	780.8	us,
'0' after	782.1	us, '1' after	782.4	us,
'0' after	783.7	us, '1' after	784	us,
'0' after	785.3	us, '1' after	797.6	us,
'0' after	798.9	us, '1' after	799.2	us,
'0' after	800.5	us, '1' after	800.8	us,
'0' after	802.1	us, '1' after	802.4	us,
'0' after	804.5	us, '1' after	816	us,
'0' after	817.3	us, '1' after	817.6	us,
'0' after	818.9	us, '1' after	819.2	us,
'0' after	821.3	us, '1' after	6806.4	us,
'0' after	6807.7	us, '1' after	6808	us,
'0' after	6809.3	us, '1' after	6809.6	us,
'0' after	6810.9	us, '1' after	6824.8	us,
'0' after	6826.1	us, '1' after	6826.4	us,
'0' after	6827.7	us, '1' after	6828	us,
'0' after	6829.3	us, '1' after	6830.4	us,
'0' after	6831.7	us, '1' after	6843.2	us,
'0' after	6844.5	us, '1' after	6844.8	us,
'0' after	6846.1	us, '1' after	6846.4	us,
'0' after	6847.7	us, '1' after	6848	us,
'0' after	6849.3	us, '1' after	6861.6	us,
'0' after	6862.9	us, '1' after	6863.2	us,
'0' after	6864.5	us, '1' after	6864.8	us,
'0' after	6866.1	us, '1' after	6866.4	us,
'0' after	6868.5	us, '1' after	6880	us,
'0' after	6881.3	us, '1' after	6881.6	us,
'0' after	6882.9	us, '1' after	6883.2	us,
'0' after	6885.3	us, '1' after	7085.6	us,
'0' after	7086.9	us, '1' after	7087.2	us,
'0' after	7088.5	us, '1' after	7088.8	us,
'0' after	7090.1	us, '1' after	7104	us,
'0' after	7105.3	us, '1' after	7105.6	us,
'0' after	7106.9	us, '1' after	7107.2	us,
'0' after	7108.5	us, '1' after	7109.6	us,
'0' after	7110.9	us, '1' after	7122.4	us,
'0' after	7123.7	us, '1' after	7124	us,
'0' after	7125.3	us, '1' after	7125.6	us,
'0' after	7126.9	us, '1' after	7127.2	us,
'0' after	7128.5	us, '1' after	7140.8	us,
'0' after	7142.1	us, '1' after	7142.4	us,
'0' after	7143.7	us, '1' after	7144	us,
'0' after	7145.3	us, '1' after	7145.6	us,
'0' after	7147.7	us, '1' after	7159.2	us,
'0' after	7160.5	us, '1' after	7160.8	us,
'0' after	7162.1	us, '1' after	7162.4	us,
'0' after	7164.5	us, '1' after	7335.2	us,
'0' after	7336.5	us, '1' after	7336.8	us,
'0' after	7338.1	us, '1' after	7338.4	us,
'0' after	7339.7	us, '1' after	7353.6	us,
'0' after	7354.9	us, '1' after	7355.2	us,
'0' after	7356.5	us, '1' after	7356.8	us,
'0' after	7358.1	us, '1' after	7359.2	us,
'0' after	7360.5	us, '1' after	7372	us,
'0' after	7373.3	us, '1' after	7373.6	us,
'0' after	7374.9	us, '1' after	7375.2	us,
'0' after	7376.5	us, '1' after	7376.8	us,
'0' after	7378.1	us, '1' after	7390.4	us,
'0' after	7391.7	us, '1' after	7392	us,
'0' after	7393.3	us, '1' after	7393.6	us,
'0' after	7394.9	us, '1' after	7395.2	us,
'0' after	7397.3	us, '1' after	7408.8	us,
'0' after	7410.1	us, '1' after	7410.4	us,
'0' after	7411.7	us, '1' after	7412	us,
'0' after	7414.1	us, '1' after	174475.2	us,
'0' after	174476.5	us, '1' after	174479.2	us,
'0' after	174481.3	us, '1' after	174494.4	us,
'0' after	174495.7	us, '1' after	174501.6	us,
'0' after	174505.3	us, '1' after	174512	us,
'0' after	174513.3	us, '1' after	174520.8	us,
'0' after	174522.1	us, '1' after	174530.4	us,
'0' after	174531.7	us, '1' after	174534.4	us,
'0' after	174538.1	us, '1' after	174548.8	us,
'0' after	174550.1	us, '1' after	174552	us,
'0' after	174553.3	us, '1' after	174553.6	us,
'0' after	174554.9	us, '1' after	174567.2	us,
'0' after	174568.5	us, '1' after	174570.4	us,
'0' after	174572.5	us, '1' after	174577.6	us,
'0' after	174578.9	us, '1' after	174585.6	us,
'0' after	174586.9	us, '1' after	174588	us,
'0' after	174589.3	us, '1' after	174604	us,
'0' after	174605.3	us, '1' after	174605.6	us,
'0' after	174608.5	us, '1' after	174608.8	us,
'0' after	174610.9	us, '1' after	174611.2	us,
'0' after	174615.7	us;




BARO_SERCLK_exp <= '0' after	2.9	us, '1' after	3.2	us,
'0' after	3.7	us, '1' after	4	us,
'0' after	4.5	us, '1' after	4.8	us,
'0' after	5.3	us, '1' after	5.6	us,
'0' after	6.1	us, '1' after	6.4	us,
'0' after	6.9	us, '1' after	7.2	us,
'0' after	7.7	us, '1' after	8	us,
'0' after	8.5	us, '1' after	8.8	us,
'0' after	9.3	us, '1' after	9.6	us,
'0' after	10.1	us, '1' after	10.4	us,
'0' after	10.9	us, '1' after	11.2	us,
'0' after	11.7	us, '1' after	12	us,
'0' after	12.5	us, '1' after	12.8	us,
'0' after	13.3	us, '1' after	13.6	us,
'0' after	14.1	us, '1' after	14.4	us,
'0' after	14.9	us, '1' after	15.2	us,
'0' after	21.3	us, '1' after	21.6	us,
'0' after	22.1	us, '1' after	22.4	us,
'0' after	22.9	us, '1' after	23.2	us,
'0' after	23.7	us, '1' after	24	us,
'0' after	24.5	us, '1' after	24.8	us,
'0' after	25.3	us, '1' after	25.6	us,
'0' after	26.1	us, '1' after	26.4	us,
'0' after	26.9	us, '1' after	27.2	us,
'0' after	27.7	us, '1' after	28	us,
'0' after	28.5	us, '1' after	28.8	us,
'0' after	29.3	us, '1' after	29.6	us,
'0' after	30.1	us, '1' after	30.4	us,
'0' after	30.9	us, '1' after	31.2	us,
'0' after	31.7	us, '1' after	32	us,
'0' after	32.5	us, '1' after	32.8	us,
'0' after	33.3	us, '1' after	33.6	us,
'0' after	39.7	us, '1' after	40	us,
'0' after	40.5	us, '1' after	40.8	us,
'0' after	41.3	us, '1' after	41.6	us,
'0' after	42.1	us, '1' after	42.4	us,
'0' after	42.9	us, '1' after	43.2	us,
'0' after	43.7	us, '1' after	44	us,
'0' after	44.5	us, '1' after	44.8	us,
'0' after	45.3	us, '1' after	45.6	us,
'0' after	46.1	us, '1' after	46.4	us,
'0' after	46.9	us, '1' after	47.2	us,
'0' after	47.7	us, '1' after	48	us,
'0' after	48.5	us, '1' after	48.8	us,
'0' after	49.3	us, '1' after	49.6	us,
'0' after	50.1	us, '1' after	50.4	us,
'0' after	50.9	us, '1' after	51.2	us,
'0' after	51.7	us, '1' after	52	us,
'0' after	58.1	us, '1' after	58.4	us,
'0' after	58.9	us, '1' after	59.2	us,
'0' after	59.7	us, '1' after	60	us,
'0' after	60.5	us, '1' after	60.8	us,
'0' after	61.3	us, '1' after	61.6	us,
'0' after	62.1	us, '1' after	62.4	us,
'0' after	62.9	us, '1' after	63.2	us,
'0' after	63.7	us, '1' after	64	us,
'0' after	64.5	us, '1' after	64.8	us,
'0' after	65.3	us, '1' after	65.6	us,
'0' after	66.1	us, '1' after	66.4	us,
'0' after	66.9	us, '1' after	67.2	us,
'0' after	67.7	us, '1' after	68	us,
'0' after	68.5	us, '1' after	68.8	us,
'0' after	69.3	us, '1' after	69.6	us,
'0' after	70.1	us, '1' after	70.4	us,
'0' after	76.5	us, '1' after	76.8	us,
'0' after	77.3	us, '1' after	77.6	us,
'0' after	78.1	us, '1' after	78.4	us,
'0' after	78.9	us, '1' after	79.2	us,
'0' after	79.7	us, '1' after	80	us,
'0' after	80.5	us, '1' after	80.8	us,
'0' after	81.3	us, '1' after	81.6	us,
'0' after	82.1	us, '1' after	82.4	us,
'0' after	82.9	us, '1' after	83.2	us,
'0' after	83.7	us, '1' after	84	us,
'0' after	84.5	us, '1' after	84.8	us,
'0' after	85.3	us, '1' after	85.6	us,
'0' after	86.1	us, '1' after	86.4	us,
'0' after	86.9	us, '1' after	87.2	us,
'0' after	87.7	us, '1' after	88	us,
'0' after	88.5	us, '1' after	88.8	us,
'0' after	94.9	us, '1' after	95.2	us,
'0' after	95.7	us, '1' after	96	us,
'0' after	96.5	us, '1' after	96.8	us,
'0' after	97.3	us, '1' after	97.6	us,
'0' after	98.1	us, '1' after	98.4	us,
'0' after	98.9	us, '1' after	99.2	us,
'0' after	99.7	us, '1' after	100	us,
'0' after	100.5	us, '1' after	100.8	us,
'0' after	101.3	us, '1' after	101.6	us,
'0' after	102.1	us, '1' after	102.4	us,
'0' after	102.9	us, '1' after	103.2	us,
'0' after	103.7	us, '1' after	104	us,
'0' after	104.5	us, '1' after	104.8	us,
'0' after	105.3	us, '1' after	105.6	us,
'0' after	106.1	us, '1' after	106.4	us,
'0' after	106.9	us, '1' after	107.2	us,
'0' after	113.3	us, '1' after	113.6	us,
'0' after	114.1	us, '1' after	114.4	us,
'0' after	114.9	us, '1' after	115.2	us,
'0' after	115.7	us, '1' after	116	us,
'0' after	116.5	us, '1' after	116.8	us,
'0' after	117.3	us, '1' after	117.6	us,
'0' after	118.1	us, '1' after	118.4	us,
'0' after	118.9	us, '1' after	119.2	us,
'0' after	119.7	us, '1' after	120	us,
'0' after	120.5	us, '1' after	120.8	us,
'0' after	121.3	us, '1' after	121.6	us,
'0' after	122.1	us, '1' after	122.4	us,
'0' after	122.9	us, '1' after	123.2	us,
'0' after	123.7	us, '1' after	124	us,
'0' after	124.5	us, '1' after	124.8	us,
'0' after	125.3	us, '1' after	125.6	us,
'0' after	131.7	us, '1' after	132	us,
'0' after	132.5	us, '1' after	132.8	us,
'0' after	133.3	us, '1' after	133.6	us,
'0' after	134.1	us, '1' after	134.4	us,
'0' after	134.9	us, '1' after	135.2	us,
'0' after	135.7	us, '1' after	136	us,
'0' after	136.5	us, '1' after	136.8	us,
'0' after	137.3	us, '1' after	137.6	us,
'0' after	138.1	us, '1' after	138.4	us,
'0' after	138.9	us, '1' after	139.2	us,
'0' after	139.7	us, '1' after	140	us,
'0' after	140.5	us, '1' after	140.8	us,
'0' after	141.3	us, '1' after	141.6	us,
'0' after	142.1	us, '1' after	142.4	us,
'0' after	142.9	us, '1' after	143.2	us,
'0' after	143.7	us, '1' after	144	us,
'0' after	166.1	us, '1' after	166.4	us,
'0' after	166.9	us, '1' after	167.2	us,
'0' after	167.7	us, '1' after	168	us,
'0' after	168.5	us, '1' after	168.8	us,
'0' after	169.3	us, '1' after	169.6	us,
'0' after	170.1	us, '1' after	170.4	us,
'0' after	170.9	us, '1' after	171.2	us,
'0' after	171.7	us, '1' after	172	us,
'0' after	172.5	us, '1' after	172.8	us,
'0' after	173.3	us, '1' after	173.6	us,
'0' after	174.1	us, '1' after	174.4	us,
'0' after	174.9	us, '1' after	175.2	us,
'0' after	175.7	us, '1' after	176	us,
'0' after	176.5	us, '1' after	176.8	us,
'0' after	177.3	us, '1' after	177.6	us,
'0' after	178.1	us, '1' after	178.4	us,
'0' after	184.5	us, '1' after	184.8	us,
'0' after	185.3	us, '1' after	185.6	us,
'0' after	186.1	us, '1' after	186.4	us,
'0' after	186.9	us, '1' after	187.2	us,
'0' after	187.7	us, '1' after	188	us,
'0' after	188.5	us, '1' after	188.8	us,
'0' after	189.3	us, '1' after	189.6	us,
'0' after	190.1	us, '1' after	190.4	us,
'0' after	190.9	us, '1' after	191.2	us,
'0' after	191.7	us, '1' after	192	us,
'0' after	192.5	us, '1' after	192.8	us,
'0' after	193.3	us, '1' after	193.6	us,
'0' after	194.1	us, '1' after	194.4	us,
'0' after	194.9	us, '1' after	195.2	us,
'0' after	195.7	us, '1' after	196	us,
'0' after	196.5	us, '1' after	196.8	us,
'0' after	202.9	us, '1' after	203.2	us,
'0' after	203.7	us, '1' after	204	us,
'0' after	204.5	us, '1' after	204.8	us,
'0' after	205.3	us, '1' after	205.6	us,
'0' after	206.1	us, '1' after	206.4	us,
'0' after	206.9	us, '1' after	207.2	us,
'0' after	207.7	us, '1' after	208	us,
'0' after	208.5	us, '1' after	208.8	us,
'0' after	209.3	us, '1' after	209.6	us,
'0' after	210.1	us, '1' after	210.4	us,
'0' after	210.9	us, '1' after	211.2	us,
'0' after	211.7	us, '1' after	212	us,
'0' after	212.5	us, '1' after	212.8	us,
'0' after	213.3	us, '1' after	213.6	us,
'0' after	214.1	us, '1' after	214.4	us,
'0' after	214.9	us, '1' after	215.2	us,
'0' after	221.3	us, '1' after	221.6	us,
'0' after	222.1	us, '1' after	222.4	us,
'0' after	222.9	us, '1' after	223.2	us,
'0' after	223.7	us, '1' after	224	us,
'0' after	224.5	us, '1' after	224.8	us,
'0' after	225.3	us, '1' after	225.6	us,
'0' after	226.1	us, '1' after	226.4	us,
'0' after	226.9	us, '1' after	227.2	us,
'0' after	227.7	us, '1' after	228	us,
'0' after	228.5	us, '1' after	228.8	us,
'0' after	229.3	us, '1' after	229.6	us,
'0' after	230.1	us, '1' after	230.4	us,
'0' after	230.9	us, '1' after	231.2	us,
'0' after	231.7	us, '1' after	232	us,
'0' after	232.5	us, '1' after	232.8	us,
'0' after	233.3	us, '1' after	233.6	us,
'0' after	239.7	us, '1' after	240	us,
'0' after	240.5	us, '1' after	240.8	us,
'0' after	241.3	us, '1' after	241.6	us,
'0' after	242.1	us, '1' after	242.4	us,
'0' after	242.9	us, '1' after	243.2	us,
'0' after	243.7	us, '1' after	244	us,
'0' after	244.5	us, '1' after	244.8	us,
'0' after	245.3	us, '1' after	245.6	us,
'0' after	246.1	us, '1' after	246.4	us,
'0' after	246.9	us, '1' after	247.2	us,
'0' after	247.7	us, '1' after	248	us,
'0' after	248.5	us, '1' after	248.8	us,
'0' after	249.3	us, '1' after	249.6	us,
'0' after	250.1	us, '1' after	250.4	us,
'0' after	250.9	us, '1' after	251.2	us,
'0' after	251.7	us, '1' after	252	us,
'0' after	742.9	us, '1' after	743.2	us,
'0' after	743.7	us, '1' after	744	us,
'0' after	744.5	us, '1' after	744.8	us,
'0' after	745.3	us, '1' after	745.6	us,
'0' after	746.1	us, '1' after	746.4	us,
'0' after	746.9	us, '1' after	747.2	us,
'0' after	747.7	us, '1' after	748	us,
'0' after	748.5	us, '1' after	748.8	us,
'0' after	749.3	us, '1' after	749.6	us,
'0' after	750.1	us, '1' after	750.4	us,
'0' after	750.9	us, '1' after	751.2	us,
'0' after	751.7	us, '1' after	752	us,
'0' after	752.5	us, '1' after	752.8	us,
'0' after	753.3	us, '1' after	753.6	us,
'0' after	754.1	us, '1' after	754.4	us,
'0' after	754.9	us, '1' after	755.2	us,
'0' after	761.3	us, '1' after	761.6	us,
'0' after	762.1	us, '1' after	762.4	us,
'0' after	762.9	us, '1' after	763.2	us,
'0' after	763.7	us, '1' after	764	us,
'0' after	764.5	us, '1' after	764.8	us,
'0' after	765.3	us, '1' after	765.6	us,
'0' after	766.1	us, '1' after	766.4	us,
'0' after	766.9	us, '1' after	767.2	us,
'0' after	767.7	us, '1' after	768	us,
'0' after	768.5	us, '1' after	768.8	us,
'0' after	769.3	us, '1' after	769.6	us,
'0' after	770.1	us, '1' after	770.4	us,
'0' after	770.9	us, '1' after	771.2	us,
'0' after	771.7	us, '1' after	772	us,
'0' after	772.5	us, '1' after	772.8	us,
'0' after	773.3	us, '1' after	773.6	us,
'0' after	779.7	us, '1' after	780	us,
'0' after	780.5	us, '1' after	780.8	us,
'0' after	781.3	us, '1' after	781.6	us,
'0' after	782.1	us, '1' after	782.4	us,
'0' after	782.9	us, '1' after	783.2	us,
'0' after	783.7	us, '1' after	784	us,
'0' after	784.5	us, '1' after	784.8	us,
'0' after	785.3	us, '1' after	785.6	us,
'0' after	786.1	us, '1' after	786.4	us,
'0' after	786.9	us, '1' after	787.2	us,
'0' after	787.7	us, '1' after	788	us,
'0' after	788.5	us, '1' after	788.8	us,
'0' after	789.3	us, '1' after	789.6	us,
'0' after	790.1	us, '1' after	790.4	us,
'0' after	790.9	us, '1' after	791.2	us,
'0' after	791.7	us, '1' after	792	us,
'0' after	798.1	us, '1' after	798.4	us,
'0' after	798.9	us, '1' after	799.2	us,
'0' after	799.7	us, '1' after	800	us,
'0' after	800.5	us, '1' after	800.8	us,
'0' after	801.3	us, '1' after	801.6	us,
'0' after	802.1	us, '1' after	802.4	us,
'0' after	802.9	us, '1' after	803.2	us,
'0' after	803.7	us, '1' after	804	us,
'0' after	804.5	us, '1' after	804.8	us,
'0' after	805.3	us, '1' after	805.6	us,
'0' after	806.1	us, '1' after	806.4	us,
'0' after	806.9	us, '1' after	807.2	us,
'0' after	807.7	us, '1' after	808	us,
'0' after	808.5	us, '1' after	808.8	us,
'0' after	809.3	us, '1' after	809.6	us,
'0' after	810.1	us, '1' after	810.4	us,
'0' after	816.5	us, '1' after	816.8	us,
'0' after	817.3	us, '1' after	817.6	us,
'0' after	818.1	us, '1' after	818.4	us,
'0' after	818.9	us, '1' after	819.2	us,
'0' after	819.7	us, '1' after	820	us,
'0' after	820.5	us, '1' after	820.8	us,
'0' after	821.3	us, '1' after	821.6	us,
'0' after	822.1	us, '1' after	822.4	us,
'0' after	822.9	us, '1' after	823.2	us,
'0' after	823.7	us, '1' after	824	us,
'0' after	824.5	us, '1' after	824.8	us,
'0' after	825.3	us, '1' after	825.6	us,
'0' after	826.1	us, '1' after	826.4	us,
'0' after	826.9	us, '1' after	827.2	us,
'0' after	827.7	us, '1' after	828	us,
'0' after	828.5	us, '1' after	828.8	us,
'0' after	6806.9	us, '1' after	6807.2	us,
'0' after	6807.7	us, '1' after	6808	us,
'0' after	6808.5	us, '1' after	6808.8	us,
'0' after	6809.3	us, '1' after	6809.6	us,
'0' after	6810.1	us, '1' after	6810.4	us,
'0' after	6810.9	us, '1' after	6811.2	us,
'0' after	6811.7	us, '1' after	6812	us,
'0' after	6812.5	us, '1' after	6812.8	us,
'0' after	6813.3	us, '1' after	6813.6	us,
'0' after	6814.1	us, '1' after	6814.4	us,
'0' after	6814.9	us, '1' after	6815.2	us,
'0' after	6815.7	us, '1' after	6816	us,
'0' after	6816.5	us, '1' after	6816.8	us,
'0' after	6817.3	us, '1' after	6817.6	us,
'0' after	6818.1	us, '1' after	6818.4	us,
'0' after	6818.9	us, '1' after	6819.2	us,
'0' after	6825.3	us, '1' after	6825.6	us,
'0' after	6826.1	us, '1' after	6826.4	us,
'0' after	6826.9	us, '1' after	6827.2	us,
'0' after	6827.7	us, '1' after	6828	us,
'0' after	6828.5	us, '1' after	6828.8	us,
'0' after	6829.3	us, '1' after	6829.6	us,
'0' after	6830.1	us, '1' after	6830.4	us,
'0' after	6830.9	us, '1' after	6831.2	us,
'0' after	6831.7	us, '1' after	6832	us,
'0' after	6832.5	us, '1' after	6832.8	us,
'0' after	6833.3	us, '1' after	6833.6	us,
'0' after	6834.1	us, '1' after	6834.4	us,
'0' after	6834.9	us, '1' after	6835.2	us,
'0' after	6835.7	us, '1' after	6836	us,
'0' after	6836.5	us, '1' after	6836.8	us,
'0' after	6837.3	us, '1' after	6837.6	us,
'0' after	6843.7	us, '1' after	6844	us,
'0' after	6844.5	us, '1' after	6844.8	us,
'0' after	6845.3	us, '1' after	6845.6	us,
'0' after	6846.1	us, '1' after	6846.4	us,
'0' after	6846.9	us, '1' after	6847.2	us,
'0' after	6847.7	us, '1' after	6848	us,
'0' after	6848.5	us, '1' after	6848.8	us,
'0' after	6849.3	us, '1' after	6849.6	us,
'0' after	6850.1	us, '1' after	6850.4	us,
'0' after	6850.9	us, '1' after	6851.2	us,
'0' after	6851.7	us, '1' after	6852	us,
'0' after	6852.5	us, '1' after	6852.8	us,
'0' after	6853.3	us, '1' after	6853.6	us,
'0' after	6854.1	us, '1' after	6854.4	us,
'0' after	6854.9	us, '1' after	6855.2	us,
'0' after	6855.7	us, '1' after	6856	us,
'0' after	6862.1	us, '1' after	6862.4	us,
'0' after	6862.9	us, '1' after	6863.2	us,
'0' after	6863.7	us, '1' after	6864	us,
'0' after	6864.5	us, '1' after	6864.8	us,
'0' after	6865.3	us, '1' after	6865.6	us,
'0' after	6866.1	us, '1' after	6866.4	us,
'0' after	6866.9	us, '1' after	6867.2	us,
'0' after	6867.7	us, '1' after	6868	us,
'0' after	6868.5	us, '1' after	6868.8	us,
'0' after	6869.3	us, '1' after	6869.6	us,
'0' after	6870.1	us, '1' after	6870.4	us,
'0' after	6870.9	us, '1' after	6871.2	us,
'0' after	6871.7	us, '1' after	6872	us,
'0' after	6872.5	us, '1' after	6872.8	us,
'0' after	6873.3	us, '1' after	6873.6	us,
'0' after	6874.1	us, '1' after	6874.4	us,
'0' after	6880.5	us, '1' after	6880.8	us,
'0' after	6881.3	us, '1' after	6881.6	us,
'0' after	6882.1	us, '1' after	6882.4	us,
'0' after	6882.9	us, '1' after	6883.2	us,
'0' after	6883.7	us, '1' after	6884	us,
'0' after	6884.5	us, '1' after	6884.8	us,
'0' after	6885.3	us, '1' after	6885.6	us,
'0' after	6886.1	us, '1' after	6886.4	us,
'0' after	6886.9	us, '1' after	6887.2	us,
'0' after	6887.7	us, '1' after	6888	us,
'0' after	6888.5	us, '1' after	6888.8	us,
'0' after	6889.3	us, '1' after	6889.6	us,
'0' after	6890.1	us, '1' after	6890.4	us,
'0' after	6890.9	us, '1' after	6891.2	us,
'0' after	6891.7	us, '1' after	6892	us,
'0' after	6892.5	us, '1' after	6892.8	us,
'0' after	7086.1	us, '1' after	7086.4	us,
'0' after	7086.9	us, '1' after	7087.2	us,
'0' after	7087.7	us, '1' after	7088	us,
'0' after	7088.5	us, '1' after	7088.8	us,
'0' after	7089.3	us, '1' after	7089.6	us,
'0' after	7090.1	us, '1' after	7090.4	us,
'0' after	7090.9	us, '1' after	7091.2	us,
'0' after	7091.7	us, '1' after	7092	us,
'0' after	7092.5	us, '1' after	7092.8	us,
'0' after	7093.3	us, '1' after	7093.6	us,
'0' after	7094.1	us, '1' after	7094.4	us,
'0' after	7094.9	us, '1' after	7095.2	us,
'0' after	7095.7	us, '1' after	7096	us,
'0' after	7096.5	us, '1' after	7096.8	us,
'0' after	7097.3	us, '1' after	7097.6	us,
'0' after	7098.1	us, '1' after	7098.4	us,
'0' after	7104.5	us, '1' after	7104.8	us,
'0' after	7105.3	us, '1' after	7105.6	us,
'0' after	7106.1	us, '1' after	7106.4	us,
'0' after	7106.9	us, '1' after	7107.2	us,
'0' after	7107.7	us, '1' after	7108	us,
'0' after	7108.5	us, '1' after	7108.8	us,
'0' after	7109.3	us, '1' after	7109.6	us,
'0' after	7110.1	us, '1' after	7110.4	us,
'0' after	7110.9	us, '1' after	7111.2	us,
'0' after	7111.7	us, '1' after	7112	us,
'0' after	7112.5	us, '1' after	7112.8	us,
'0' after	7113.3	us, '1' after	7113.6	us,
'0' after	7114.1	us, '1' after	7114.4	us,
'0' after	7114.9	us, '1' after	7115.2	us,
'0' after	7115.7	us, '1' after	7116	us,
'0' after	7116.5	us, '1' after	7116.8	us,
'0' after	7122.9	us, '1' after	7123.2	us,
'0' after	7123.7	us, '1' after	7124	us,
'0' after	7124.5	us, '1' after	7124.8	us,
'0' after	7125.3	us, '1' after	7125.6	us,
'0' after	7126.1	us, '1' after	7126.4	us,
'0' after	7126.9	us, '1' after	7127.2	us,
'0' after	7127.7	us, '1' after	7128	us,
'0' after	7128.5	us, '1' after	7128.8	us,
'0' after	7129.3	us, '1' after	7129.6	us,
'0' after	7130.1	us, '1' after	7130.4	us,
'0' after	7130.9	us, '1' after	7131.2	us,
'0' after	7131.7	us, '1' after	7132	us,
'0' after	7132.5	us, '1' after	7132.8	us,
'0' after	7133.3	us, '1' after	7133.6	us,
'0' after	7134.1	us, '1' after	7134.4	us,
'0' after	7134.9	us, '1' after	7135.2	us,
'0' after	7141.3	us, '1' after	7141.6	us,
'0' after	7142.1	us, '1' after	7142.4	us,
'0' after	7142.9	us, '1' after	7143.2	us,
'0' after	7143.7	us, '1' after	7144	us,
'0' after	7144.5	us, '1' after	7144.8	us,
'0' after	7145.3	us, '1' after	7145.6	us,
'0' after	7146.1	us, '1' after	7146.4	us,
'0' after	7146.9	us, '1' after	7147.2	us,
'0' after	7147.7	us, '1' after	7148	us,
'0' after	7148.5	us, '1' after	7148.8	us,
'0' after	7149.3	us, '1' after	7149.6	us,
'0' after	7150.1	us, '1' after	7150.4	us,
'0' after	7150.9	us, '1' after	7151.2	us,
'0' after	7151.7	us, '1' after	7152	us,
'0' after	7152.5	us, '1' after	7152.8	us,
'0' after	7153.3	us, '1' after	7153.6	us,
'0' after	7159.7	us, '1' after	7160	us,
'0' after	7160.5	us, '1' after	7160.8	us,
'0' after	7161.3	us, '1' after	7161.6	us,
'0' after	7162.1	us, '1' after	7162.4	us,
'0' after	7162.9	us, '1' after	7163.2	us,
'0' after	7163.7	us, '1' after	7164	us,
'0' after	7164.5	us, '1' after	7164.8	us,
'0' after	7165.3	us, '1' after	7165.6	us,
'0' after	7166.1	us, '1' after	7166.4	us,
'0' after	7166.9	us, '1' after	7167.2	us,
'0' after	7167.7	us, '1' after	7168	us,
'0' after	7168.5	us, '1' after	7168.8	us,
'0' after	7169.3	us, '1' after	7169.6	us,
'0' after	7170.1	us, '1' after	7170.4	us,
'0' after	7170.9	us, '1' after	7171.2	us,
'0' after	7171.7	us, '1' after	7172	us,
'0' after	7335.7	us, '1' after	7336	us,
'0' after	7336.5	us, '1' after	7336.8	us,
'0' after	7337.3	us, '1' after	7337.6	us,
'0' after	7338.1	us, '1' after	7338.4	us,
'0' after	7338.9	us, '1' after	7339.2	us,
'0' after	7339.7	us, '1' after	7340	us,
'0' after	7340.5	us, '1' after	7340.8	us,
'0' after	7341.3	us, '1' after	7341.6	us,
'0' after	7342.1	us, '1' after	7342.4	us,
'0' after	7342.9	us, '1' after	7343.2	us,
'0' after	7343.7	us, '1' after	7344	us,
'0' after	7344.5	us, '1' after	7344.8	us,
'0' after	7345.3	us, '1' after	7345.6	us,
'0' after	7346.1	us, '1' after	7346.4	us,
'0' after	7346.9	us, '1' after	7347.2	us,
'0' after	7347.7	us, '1' after	7348	us,
'0' after	7354.1	us, '1' after	7354.4	us,
'0' after	7354.9	us, '1' after	7355.2	us,
'0' after	7355.7	us, '1' after	7356	us,
'0' after	7356.5	us, '1' after	7356.8	us,
'0' after	7357.3	us, '1' after	7357.6	us,
'0' after	7358.1	us, '1' after	7358.4	us,
'0' after	7358.9	us, '1' after	7359.2	us,
'0' after	7359.7	us, '1' after	7360	us,
'0' after	7360.5	us, '1' after	7360.8	us,
'0' after	7361.3	us, '1' after	7361.6	us,
'0' after	7362.1	us, '1' after	7362.4	us,
'0' after	7362.9	us, '1' after	7363.2	us,
'0' after	7363.7	us, '1' after	7364	us,
'0' after	7364.5	us, '1' after	7364.8	us,
'0' after	7365.3	us, '1' after	7365.6	us,
'0' after	7366.1	us, '1' after	7366.4	us,
'0' after	7372.5	us, '1' after	7372.8	us,
'0' after	7373.3	us, '1' after	7373.6	us,
'0' after	7374.1	us, '1' after	7374.4	us,
'0' after	7374.9	us, '1' after	7375.2	us,
'0' after	7375.7	us, '1' after	7376	us,
'0' after	7376.5	us, '1' after	7376.8	us,
'0' after	7377.3	us, '1' after	7377.6	us,
'0' after	7378.1	us, '1' after	7378.4	us,
'0' after	7378.9	us, '1' after	7379.2	us,
'0' after	7379.7	us, '1' after	7380	us,
'0' after	7380.5	us, '1' after	7380.8	us,
'0' after	7381.3	us, '1' after	7381.6	us,
'0' after	7382.1	us, '1' after	7382.4	us,
'0' after	7382.9	us, '1' after	7383.2	us,
'0' after	7383.7	us, '1' after	7384	us,
'0' after	7384.5	us, '1' after	7384.8	us,
'0' after	7390.9	us, '1' after	7391.2	us,
'0' after	7391.7	us, '1' after	7392	us,
'0' after	7392.5	us, '1' after	7392.8	us,
'0' after	7393.3	us, '1' after	7393.6	us,
'0' after	7394.1	us, '1' after	7394.4	us,
'0' after	7394.9	us, '1' after	7395.2	us,
'0' after	7395.7	us, '1' after	7396	us,
'0' after	7396.5	us, '1' after	7396.8	us,
'0' after	7397.3	us, '1' after	7397.6	us,
'0' after	7398.1	us, '1' after	7398.4	us,
'0' after	7398.9	us, '1' after	7399.2	us,
'0' after	7399.7	us, '1' after	7400	us,
'0' after	7400.5	us, '1' after	7400.8	us,
'0' after	7401.3	us, '1' after	7401.6	us,
'0' after	7402.1	us, '1' after	7402.4	us,
'0' after	7402.9	us, '1' after	7403.2	us,
'0' after	7409.3	us, '1' after	7409.6	us,
'0' after	7410.1	us, '1' after	7410.4	us,
'0' after	7410.9	us, '1' after	7411.2	us,
'0' after	7411.7	us, '1' after	7412	us,
'0' after	7412.5	us, '1' after	7412.8	us,
'0' after	7413.3	us, '1' after	7413.6	us,
'0' after	7414.1	us, '1' after	7414.4	us,
'0' after	7414.9	us, '1' after	7415.2	us,
'0' after	7415.7	us, '1' after	7416	us,
'0' after	7416.5	us, '1' after	7416.8	us,
'0' after	7417.3	us, '1' after	7417.6	us,
'0' after	7418.1	us, '1' after	7418.4	us,
'0' after	7418.9	us, '1' after	7419.2	us,
'0' after	7419.7	us, '1' after	7420	us,
'0' after	7420.5	us, '1' after	7420.8	us,
'0' after	7421.3	us, '1' after	7421.6	us,
'0' after	174474.1	us, '1' after	174474.4	us,
'0' after	174474.9	us, '1' after	174475.2	us,
'0' after	174475.7	us, '1' after	174476	us,
'0' after	174476.5	us, '1' after	174476.8	us,
'0' after	174477.3	us, '1' after	174477.6	us,
'0' after	174478.1	us, '1' after	174478.4	us,
'0' after	174478.9	us, '1' after	174479.2	us,
'0' after	174479.7	us, '1' after	174480	us,
'0' after	174480.5	us, '1' after	174480.8	us,
'0' after	174481.3	us, '1' after	174481.6	us,
'0' after	174482.1	us, '1' after	174482.4	us,
'0' after	174482.9	us, '1' after	174483.2	us,
'0' after	174483.7	us, '1' after	174484	us,
'0' after	174484.5	us, '1' after	174484.8	us,
'0' after	174485.3	us, '1' after	174485.6	us,
'0' after	174486.1	us, '1' after	174486.4	us,
'0' after	174492.5	us, '1' after	174492.8	us,
'0' after	174493.3	us, '1' after	174493.6	us,
'0' after	174494.1	us, '1' after	174494.4	us,
'0' after	174494.9	us, '1' after	174495.2	us,
'0' after	174495.7	us, '1' after	174496	us,
'0' after	174496.5	us, '1' after	174496.8	us,
'0' after	174497.3	us, '1' after	174497.6	us,
'0' after	174498.1	us, '1' after	174498.4	us,
'0' after	174498.9	us, '1' after	174499.2	us,
'0' after	174499.7	us, '1' after	174500	us,
'0' after	174500.5	us, '1' after	174500.8	us,
'0' after	174501.3	us, '1' after	174501.6	us,
'0' after	174502.1	us, '1' after	174502.4	us,
'0' after	174502.9	us, '1' after	174503.2	us,
'0' after	174503.7	us, '1' after	174504	us,
'0' after	174504.5	us, '1' after	174504.8	us,
'0' after	174510.9	us, '1' after	174511.2	us,
'0' after	174511.7	us, '1' after	174512	us,
'0' after	174512.5	us, '1' after	174512.8	us,
'0' after	174513.3	us, '1' after	174513.6	us,
'0' after	174514.1	us, '1' after	174514.4	us,
'0' after	174514.9	us, '1' after	174515.2	us,
'0' after	174515.7	us, '1' after	174516	us,
'0' after	174516.5	us, '1' after	174516.8	us,
'0' after	174517.3	us, '1' after	174517.6	us,
'0' after	174518.1	us, '1' after	174518.4	us,
'0' after	174518.9	us, '1' after	174519.2	us,
'0' after	174519.7	us, '1' after	174520	us,
'0' after	174520.5	us, '1' after	174520.8	us,
'0' after	174521.3	us, '1' after	174521.6	us,
'0' after	174522.1	us, '1' after	174522.4	us,
'0' after	174522.9	us, '1' after	174523.2	us,
'0' after	174529.3	us, '1' after	174529.6	us,
'0' after	174530.1	us, '1' after	174530.4	us,
'0' after	174530.9	us, '1' after	174531.2	us,
'0' after	174531.7	us, '1' after	174532	us,
'0' after	174532.5	us, '1' after	174532.8	us,
'0' after	174533.3	us, '1' after	174533.6	us,
'0' after	174534.1	us, '1' after	174534.4	us,
'0' after	174534.9	us, '1' after	174535.2	us,
'0' after	174535.7	us, '1' after	174536	us,
'0' after	174536.5	us, '1' after	174536.8	us,
'0' after	174537.3	us, '1' after	174537.6	us,
'0' after	174538.1	us, '1' after	174538.4	us,
'0' after	174538.9	us, '1' after	174539.2	us,
'0' after	174539.7	us, '1' after	174540	us,
'0' after	174540.5	us, '1' after	174540.8	us,
'0' after	174541.3	us, '1' after	174541.6	us,
'0' after	174547.7	us, '1' after	174548	us,
'0' after	174548.5	us, '1' after	174548.8	us,
'0' after	174549.3	us, '1' after	174549.6	us,
'0' after	174550.1	us, '1' after	174550.4	us,
'0' after	174550.9	us, '1' after	174551.2	us,
'0' after	174551.7	us, '1' after	174552	us,
'0' after	174552.5	us, '1' after	174552.8	us,
'0' after	174553.3	us, '1' after	174553.6	us,
'0' after	174554.1	us, '1' after	174554.4	us,
'0' after	174554.9	us, '1' after	174555.2	us,
'0' after	174555.7	us, '1' after	174556	us,
'0' after	174556.5	us, '1' after	174556.8	us,
'0' after	174557.3	us, '1' after	174557.6	us,
'0' after	174558.1	us, '1' after	174558.4	us,
'0' after	174558.9	us, '1' after	174559.2	us,
'0' after	174559.7	us, '1' after	174560	us,
'0' after	174566.1	us, '1' after	174566.4	us,
'0' after	174566.9	us, '1' after	174567.2	us,
'0' after	174567.7	us, '1' after	174568	us,
'0' after	174568.5	us, '1' after	174568.8	us,
'0' after	174569.3	us, '1' after	174569.6	us,
'0' after	174570.1	us, '1' after	174570.4	us,
'0' after	174570.9	us, '1' after	174571.2	us,
'0' after	174571.7	us, '1' after	174572	us,
'0' after	174572.5	us, '1' after	174572.8	us,
'0' after	174573.3	us, '1' after	174573.6	us,
'0' after	174574.1	us, '1' after	174574.4	us,
'0' after	174574.9	us, '1' after	174575.2	us,
'0' after	174575.7	us, '1' after	174576	us,
'0' after	174576.5	us, '1' after	174576.8	us,
'0' after	174577.3	us, '1' after	174577.6	us,
'0' after	174578.1	us, '1' after	174578.4	us,
'0' after	174584.5	us, '1' after	174584.8	us,
'0' after	174585.3	us, '1' after	174585.6	us,
'0' after	174586.1	us, '1' after	174586.4	us,
'0' after	174586.9	us, '1' after	174587.2	us,
'0' after	174587.7	us, '1' after	174588	us,
'0' after	174588.5	us, '1' after	174588.8	us,
'0' after	174589.3	us, '1' after	174589.6	us,
'0' after	174590.1	us, '1' after	174590.4	us,
'0' after	174590.9	us, '1' after	174591.2	us,
'0' after	174591.7	us, '1' after	174592	us,
'0' after	174592.5	us, '1' after	174592.8	us,
'0' after	174593.3	us, '1' after	174593.6	us,
'0' after	174594.1	us, '1' after	174594.4	us,
'0' after	174594.9	us, '1' after	174595.2	us,
'0' after	174595.7	us, '1' after	174596	us,
'0' after	174596.5	us, '1' after	174596.8	us,
'0' after	174602.9	us, '1' after	174603.2	us,
'0' after	174603.7	us, '1' after	174604	us,
'0' after	174604.5	us, '1' after	174604.8	us,
'0' after	174605.3	us, '1' after	174605.6	us,
'0' after	174606.1	us, '1' after	174606.4	us,
'0' after	174606.9	us, '1' after	174607.2	us,
'0' after	174607.7	us, '1' after	174608	us,
'0' after	174608.5	us, '1' after	174608.8	us,
'0' after	174609.3	us, '1' after	174609.6	us,
'0' after	174610.1	us, '1' after	174610.4	us,
'0' after	174610.9	us, '1' after	174611.2	us,
'0' after	174611.7	us, '1' after	174612	us,
'0' after	174612.5	us, '1' after	174612.8	us,
'0' after	174613.3	us, '1' after	174613.6	us,
'0' after	174614.1	us, '1' after	174614.4	us,
'0' after	174614.9	us, '1' after	174615.2	us;




baro_CSN_exp <= 	'1' AFTER 0 US,			
'0' after	2.1	us, '1' after	16.5	us,
'0' after	20.5	us, '1' after	34.9	us,
'0' after	38.9	us, '1' after	53.3	us,
'0' after	57.3	us, '1' after	71.7	us,
'0' after	75.7	us, '1' after	90.1	us,
'0' after	94.1	us, '1' after	108.5	us,
'0' after	112.5	us, '1' after	126.9	us,
'0' after	130.9	us, '1' after	145.3	us,
'0' after	165.3	us, '1' after	179.7	us,
'0' after	183.7	us, '1' after	198.1	us,
'0' after	202.1	us, '1' after	216.5	us,
'0' after	220.5	us, '1' after	234.9	us,
'0' after	238.9	us, '1' after	253.3	us,
'0' after	742.1	us, '1' after	756.5	us,
'0' after	760.5	us, '1' after	774.9	us,
'0' after	778.9	us, '1' after	793.3	us,
'0' after	797.3	us, '1' after	811.7	us,
'0' after	815.7	us, '1' after	830.1	us,
'0' after	174473.5	us, '1' after	147487.7	us,
'0' after	174491.9	us, '1' after	174506.1	us,
'0' after	174510.3	us, '1' after	174524.5	us,
'0' after	174528.5	us, '1' after	174542.9	us,
'0' after	174546.9	us, '1' after	174561.3	us,
'0' after	174565.5	us, '1' after	174579.7	us,
'0' after	174583.9	us, '1' after	174598.1	us,
'0' after	174602.3	us, '1' after	174616.1	us;


--Comparator

end architecture testbench;

